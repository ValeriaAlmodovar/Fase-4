//==============================================================
//  Second Operand Handler
//==============================================================
module SOH (
    input  wire [31:0] R,          // rs2 value
    input  wire [12:0] imm13,      // immediate for ALU/LD/ST
    input  wire [21:0] imm22,      // immediate for sethi / branches
    input  wire [3:0]  S,          // selector
    output reg  [31:0] N
);

always @(*) begin
    case (S)

        //===============================
        // 0000 : Use R (default)
        //===============================
        4'b0000: N = R;

        //===============================
        // 0001 : Imm13 sign-extended
        //===============================
        4'b0001: N = {{19{imm13[12]}}, imm13};

        //===============================
        // 0010 : SETHI → imm22 << 10
        //===============================
        4'b0010: N = {imm22, 10'b0};

        //===============================
        // 0011 : Branch displacement
        // disp22 << 2, sign-extended
        //===============================
        4'b0011: N = {{8{imm22[21]}}, imm22, 2'b00};

        //===============================
        // 0100 : Shift by R[4:0]
        //===============================
        4'b0100: N = {27'b0, R[4:0]};

        //===============================
        // 0101 : Shift by imm13[4:0]
        //===============================
        4'b0101: N = {27'b0, imm13[4:0]};

        //===============================
        // DEFAULT
        //===============================
        default: N = R;
    endcase
end

endmodule
