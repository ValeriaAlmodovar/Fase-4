//==============================================================
//  ALU de 32 bits 
//==============================================================
module ALU
(
    input  wire [31:0] A, B,      // Entradas de 32 bits
    input  wire        Ci,        // Carry-in 
    input  wire [3:0]  ALU_OP,    // Código reducido desde la CU

    output reg  [31:0] ALU_OUT,   // Resultado
    output reg         Z_EX,      // Zero flag
    output reg         N_EX,      // Negative flag
    output reg         C_EX,      // Carry flag
    output reg         V_EX       // Overflow flag
);

    // Resultado extendido (para detectar carry/borrow)
    reg [32:0] Result;

    // Ejecuta este bloque cada vez que cualquier entrada cambie
    always @* begin

        // Reinicialización de salidas
        ALU_OUT = 32'b0;
        Z_EX    = 1'b0;
        N_EX    = 1'b0;
        C_EX    = 1'b0;
        V_EX    = 1'b0;
        Result  = 33'b0;

        case (ALU_OP)

            //==================================================
            // 0000 : ADD   (SPARC op3 = 000000)
            //  rd ← rs1 + op2
            //==================================================
            4'b0000: begin
                Result  = {1'b0, A} + {1'b0, B};
                ALU_OUT = Result[31:0];
                C_EX    = Result[32];
                V_EX    = (~(A[31] ^ B[31])) & (A[31] ^ ALU_OUT[31]);
            end

            //==================================================
            // 0001 : addcc (SPARC op3 = 010000)
            //  rd ← rs1 + op2   
            //==================================================
            4'b0001: begin
                Result  = {1'b0, A} + {1'b0, B};
                ALU_OUT = Result[31:0];
                C_EX    = Result[32];
                V_EX    = (~(A[31] ^ B[31])) & (A[31] ^ ALU_OUT[31]);
            end

            //==================================================
            // 0010 : SUB   (SPARC op3 = 000100)
            //  rd ← rs1 - op2
            //==================================================
            4'b0010: begin
                Result  = {1'b0, A} + {1'b0, ~B} + 33'b1;  // A - B
                ALU_OUT = Result[31:0];
                C_EX    = Result[32];
                V_EX    = (A[31] ^ B[31]) & (A[31] ^ ALU_OUT[31]);
            end

            //==================================================
            // 0011 : subcc (SPARC op3 = 010100)
            //  rd ← rs1 - op2   
            //==================================================
            4'b0011: begin
                Result  = {1'b0, A} + {1'b0, ~B} + 33'b1;
                ALU_OUT = Result[31:0];
                C_EX    = Result[32];
                V_EX    = (A[31] ^ B[31]) & (A[31] ^ ALU_OUT[31]);
            end

            //==================================================
            // 0100 : AND   (SPARC op3 = 000001)
            //  rd ← rs1 & op2
            //==================================================
            4'b0100: begin
                ALU_OUT = A & B;
            end

            //==================================================
            // 0101 : OR    (SPARC op3 = 000010)
            //  rd ← rs1 | op2
            //==================================================
            4'b0101: begin
                ALU_OUT = A | B;
            end

            //==================================================
            // 0110 : XOR   (SPARC op3 = 000011)
            //  rd ← rs1 ^ op2
            //==================================================
            4'b0110: begin
                ALU_OUT = A ^ B;
            end

            //==================================================
            // 0111 : XNOR  (SPARC op3 = 000111)
            //  rd ← ~(rs1 ^ op2)
            //==================================================
            4'b0111: begin
                ALU_OUT = ~(A ^ B);
            end

            //==================================================
            // 1000 : ANDN  (SPARC op3 = 000101)
            //  rd ← rs1 & ~op2
            //==================================================
            4'b1000: begin
                ALU_OUT = A & ~B;
            end

            //==================================================
            // 1001 : ORN   (SPARC op3 = 000110)
            //  rd ← rs1 | ~op2
            //==================================================
            4'b1001: begin
                ALU_OUT = A | ~B;
            end

            //==================================================
            // 1010 : SLL   (SPARC op3 = 100101)
            //  rd ← rs1 << op2[4:0]
            //==================================================
            4'b1010: begin
                ALU_OUT = A << B[4:0];
            end

            //==================================================
            // 1011 : SRL   (SPARC op3 = 100110)
            //  rd ← rs1 >> op2[4:0]
            //==================================================
            4'b1011: begin
                ALU_OUT = A >> B[4:0];
            end

            //==================================================
            // 1100 : SRA   (SPARC op3 = 100111)
            //  rd ← rs1 >>> op2[4:0]  (sign-extend)
            //==================================================
            4'b1100: begin
                ALU_OUT = $signed(A) >>> B[4:0];
            end

            //==================================================
            // 1101 : PASS B (para SETHI)
            //  rd ← imm22 << 10
            //==================================================
            4'b1101: begin
                ALU_OUT = B;
            end

            //==================================================
            // 1110 : ADDX (ADD with carry)
            //  rd ← rs1 + op2 + Ci
            //==================================================
            4'b1110: begin
                Result  = {1'b0, A} + {1'b0, B} + {32'b0, Ci};
                ALU_OUT = Result[31:0];
                C_EX    = Result[32];
                V_EX    = (~(A[31] ^ B[31])) & (A[31] ^ ALU_OUT[31]);
            end

            //==================================================
            // 1111 : SUBX (SUB with carry/borrow)
            //  rd ← rs1 - op2 - Ci
            //==================================================
            4'b1111: begin
                Result  = {1'b0, A} + {1'b0, ~B} + {32'b0, Ci};
                ALU_OUT = Result[31:0];
                C_EX    = Result[32];
                V_EX    = (A[31] ^ B[31]) & (A[31] ^ ALU_OUT[31]);
            end

            //==================================================
            // DEFAULT
            //==================================================
            default: begin
                ALU_OUT = 32'b0;
            end
        endcase

        //==================================================
        // FLAGS siempre producidos
        // REG_CC decide si guardarlos (CC_WE)
        //==================================================
        Z_EX = (ALU_OUT == 32'b0);
        N_EX = ALU_OUT[31];
    end

endmodule
