//==============================================================
//  register_zero
//==============================================================

module register_zero (
    output wire [31:0] Q
);

assign Q = 32'b0;

endmodule
